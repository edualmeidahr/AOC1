library verilog;
use verilog.vl_types.all;
entity Register_Bank_vlg_vec_tst is
end Register_Bank_vlg_vec_tst;
